
`default_nettype none
 `define USE_PACOBLAZE
module 
picoblaze_template
#(
parameter clk_freq_in_hz = 50000000 //50MHz clock
) (
				output reg[7:0] led,
				input clk,
				input [7:0] input_data1,
        input [7:0] input_data2,
        input [7:0] input_data3,
        input [7:0] input_data4,
        input interrupt_signal,
			  output wire [23:0] sseg,
				output reg LED0
			     );


  
//--
//------------------------------------------------------------------------------------
//--
//-- Signals used to connect KCPSM3 to program ROM and I/O logic
//--

wire[9:0]  address;
wire[17:0]  instruction;
wire[7:0]  port_id;
wire[7:0]  out_port;
reg[7:0]  in_port;
wire  write_strobe;
wire  read_strobe;
reg  interrupt;
wire  interrupt_ack;
wire  kcpsm3_reset;

//--
//-- Signals used to generate interrupt (not used in lab)
//--
// reg[26:0] int_count;
// reg event_1hz;

//-- Signals for LCD operation
//--
//--

reg        lcd_rw_control;
reg[7:0]   lcd_output_data;
pacoblaze3 led_8seg_kcpsm //pacoblaze module
(
                  .address(address),
               .instruction(instruction),
                   .port_id(port_id),
              .write_strobe(write_strobe),
                  .out_port(out_port),
               .read_strobe(read_strobe),
                   .in_port(in_port),
                 .interrupt(interrupt),
             .interrupt_ack(interrupt_ack),
                     .reset(kcpsm3_reset),
                       .clk(clk));

 wire [19:0] raw_instruction;
	
	pacoblaze_instruction_memory 
	pacoblaze_instruction_memory_inst(
     	.addr(address),
	    .outdata(raw_instruction)
	);
	
	always @ (posedge clk)
	begin
	      instruction <= raw_instruction[17:0];
	end

    assign kcpsm3_reset = 0;                       
  
//  ----------------------------------------------------------------------------------------------------------------------------------
//  -- Interrupt 
//  ----------------------------------------------------------------------------------------------------------------------------------
//  --
//  --
//  -- Interrupt is used to provide a 1 second time reference.
//  --
//  --
//  -- A simple binary counter is used to divide the 50MHz system clock and provide interrupt pulses.
//  --


// Note that because we are using clock enable we DO NOT need to synchronize with clk

//   always @ (posedge clk)
//   begin
//       //--divide 50MHz by 50,000,000 to form 1Hz pulses
//       if (int_count==(clk_freq_in_hz-1)) //clock enable
//       begin
//           int_count <= 0;
//           event_1hz <= 1;
//       end else
//       begin
//           int_count <= int_count + 1;
//           event_1hz <= 0;
//       end
//  end

//Don't need, this was included in original template code, basic interrupt signal handling

//  always @ (posedge clk or posedge interrupt_ack)  //FF with clock "clk" and reset "interrupt_ack"
//  begin
//       if (interrupt_ack) //if we get reset, reset interrupt in order to wait for next clock.
//             interrupt <= 0;
//       else
// 		begin 
// 		      if (event_1hz)   //clock enable
//       		      interrupt <= 1;
//           		else
// 		            interrupt <= interrupt;
//       end
//  end


//Interrupt based on signal from top module simple_ipod_solution.v
always @ (posedge clk or posedge interrupt_ack)
begin
    if (interrupt_ack) //if interrupt reset, go to 0
        interrupt <= 0;
    else
        interrupt <= interrupt_signal; //send interrupt signal
end

//  --
//  ----------------------------------------------------------------------------------------------------------------------------------
//  -- KCPSM3 input ports 
//  ----------------------------------------------------------------------------------------------------------------------------------
//  --
//  --
//  -- The inputs connect via a pipelined multiplexer
//  --

 always @ (posedge clk)
 begin
    case (port_id[7:0]) //Input ports, input_data sent in three ports (only one actual input port, so must mux them together)
        8'h0:    in_port <= input_data1;
        8'h1:    in_port <= input_data2;
        8'h2:    in_port <= input_data3;
        8'h3:    in_port <= input_data4;
        default: in_port <= 8'bx;
    endcase
end
   
//
//  --
//  ----------------------------------------------------------------------------------------------------------------------------------
//  -- KCPSM3 output ports 
//  ----------------------------------------------------------------------------------------------------------------------------------
//  --
//  -- adding the output registers to the processor
//  --
//   
  always @ (posedge clk)
  begin

        //port 80 hex 
        if (write_strobe & port_id[7])  //LEDR[9:2] output port
          led <= out_port;

        //port 40 hex 
        if (write_strobe & port_id[6])  //clock enable 
          sseg[7:0] <= out_port;
			      
		  //port 20 hex 
		  if (write_strobe & port_id[5])  //clock enable 
          sseg[15:8] <= out_port;
			      
		  //port 10 hex 			
        if (write_strobe & port_id[4])  //clock enable 
          sseg[23:16] <= out_port;
			 
			 
		  if (write_strobe & port_id[0]) //LED0 output port
          LED0 <= out_port;
				
			      
  end

endmodule
